yyy line ttt hhh kkk
test