this file has   multiple spaces between words
spaces at the end of a line     
and  	tabs between	some 	words

it 	also has an empty line
  	 
and a line with just whitespace
