if (a /=letterB and letterB<= c and c >=d) then
b := a;
b:=a**a;
d <=letterB;
e<= a& letterB;
f <= (others=> '0');
end if;
