signal a,letterB,c,d : std_logic ;
if ( a = letterB+c-d or letterB*letterB = c or a > c) then
end if;
