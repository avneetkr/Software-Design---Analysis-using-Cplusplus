CLK'EVENT and CLK = '1'
aBit = '0' and vector ' length
