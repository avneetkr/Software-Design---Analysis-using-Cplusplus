x"00101AB010" X"01FFF0111" "0101000"
"011000" O"01237"
