CLK'EVENT
vector ' length
