CLK'EVENT
vector ' length
a=1;