signal a,letterB,c,d : std_logic(3 downto 1) ;
if ( a = letterB+c-d or letterB*letterB = c or a > c) then
end if;
