'0' '1'
'-' 'Z'
