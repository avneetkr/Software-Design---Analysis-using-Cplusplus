-- a plain comment
  --comment with tab in front
      --comment with whitespace at the end        
--comment with VHDL code inside y <= a * b;
  y <= a *b;    --comment
y <= a * b;--comment right after code
--comment with comment -- symbol inside -- --

