this file has only a single space between words
and no spaces at the end of any
line
