--comment
-- another comment
