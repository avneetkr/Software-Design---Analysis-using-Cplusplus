"00101010" "010111"
